interface Ifc_;
endinterface
